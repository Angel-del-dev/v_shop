module structs


pub struct Product{
	pub mut: 
		name string
		price f64 // float64
}